
module CPU (
	clk_clk,
	led_export);	

	input		clk_clk;
	output	[1:0]	led_export;
endmodule
