module top_control ( 
input  CLOCK_50,              // 50 MHz Clock ref
input  ADC_SDAT,              // SPI ADC MISO
output ADC_CS_N,              // SPI ADC nCS
output ADC_SADDR,             // SPI ADC MOSI
output ADC_SCLK,              // SPI ADC SCK
output GPIO_00,               // PID out PWM
output [7:0] LED
);




//////-----ADC-SPI-----//////
wire ClkDev;
wire [7:0] in_adc_chanel_read = 8'b0;         // (default) IN0
wire o_RX_DV;
wire o_TX_Ready;
wire [7:0] adc_RX_Byte;

reg [7:0] count_byte  = 0;
reg [7:0] rx_byte_MSB = 0;
reg [7:0] rx_byte_LSB = 0;

assign ADC_CS_N = 1'b0;
clock_divider #(.M(4)) (.clock_out(ClkDev), .clk_in(CLOCK_50));

spi_master
#(.SPI_MODE(0), .CLKS_PER_HALF_BIT(4))
  (
   // Control/Data Signals,
   .i_Rst_L(1'b1),                          // FPGA Reset
   .i_Clk(CLOCK_50),                        // FPGA Clock
   
   // TX (MOSI) Signals
   .i_TX_Byte(in_adc_chanel_read),          // Byte to transmit on MOSI
   .i_TX_DV(ClkDev),                        // Data Valid Pulse with i_TX_Byte
   .o_TX_Ready(o_TX_Ready),                 // Transmit Ready for next byte
   
   // RX (MISO) Signals
   .o_RX_DV(o_RX_DV),                       // Data Valid pulse (1 clock cycle)
   .o_RX_Byte(adc_RX_Byte),                 // Byte received on MISO

   // SPI Interface
   .o_SPI_Clk(ADC_SCLK),
   .i_SPI_MISO(ADC_SDAT),
   .o_SPI_MOSI(ADC_SADDR)
   );

/// --- RX MSB and LSB byte --- ///
always @(posedge ADC_SCLK)
begin
count_byte = count_byte + 1;
	if (count_byte == 1)
	begin
		rx_byte_MSB <= adc_RX_Byte;
	end
		if (count_byte == 2)
		begin
			rx_byte_LSB <= adc_RX_Byte;
			count_byte = 0;
		end
end

wire [7:0] w_rx_byte_MSB;
wire [7:0] W_rx_byte_LSB;

assign w_rx_byte_MSB = rx_byte_MSB;
assign w_rx_byte_LSB = rx_byte_LSB;

reg  [11:0] ADC_Data;
wire [11:0] w_ADC_DAta;

assign w_ADC_DAta = ADC_Data;

//// --- function calc ADC data 12-bit --- ////
function [11:0] temp_ADC_data (input [7:0] MSB, LSB);
temp_ADC_data = {MSB,LSB};   // or ((MSB<<8)|LSB);
endfunction 

/// --- 12-bit data ADC --- ///
always @(posedge CLOCK_50)
begin
	ADC_Data <= temp_ADC_data(w_rx_byte_MSB,w_rx_byte_LSB);
end

//////----PWM-OUT----///////
PWM_PID #(.DataTopValue(32767), .DataWidth(15)) (  
.PWM_outP(GPIO_00), 
.data(w_ADC_DAta), 
.clk_in(CLOCK_50),
.enable(1'b1),
.reset(1'b0));

assign LED[0] = GPIO_00; // real PWM out LED indicate

endmodule 